------------------------------------------------------------------------------
-- Taken from the documentation for GHDL.                                    |
-- See https://github.com/gritbub/learning/blob/master/fpga/vhdl/Sources.md  |
--    for license info.                                                      |
------------------------------------------------------------------------------


entity adder is
   -- i0, i1, and the carry-in ci are inputs of the adder.
   -- s is the sum output, co is the carry-out.
   port ( i0, i1, ci : in bit; s, co : out bit );
end adder;

architecture rt1 of adder is
begin
   -- This full-adder architecture contains two concurrent assignments.
   -- Compute the sum:
   s <= i0 xor i1 xor ci;
   -- Compute the carry.
   co <= (i0 and i1) or (i0 and ci) or (i1 and ci);
end rt1;

